import params_pkg::*;

module directory_controller (
    input logic aclk,
    input logic arst_n,
);

endmodule : directory_controller
